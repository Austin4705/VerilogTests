module pls(input a, output b);
        not (a, b);
endmodule